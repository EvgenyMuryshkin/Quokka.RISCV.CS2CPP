`default_nettype none

module RVTest (
	input clk,
	input resetn,
	output         o_mem_valid,
	output         o_mem_instr,

	output  [31:0] 	o_mem_addr,
	output  [31:0] 	o_mem_wdata,
	output  [ 3:0] 	o_mem_wstrb,
	output 			o_dbg_mem_valid,
	output [31:0] 	o_dbg_mem_rdata,
	output [31:0] 	o_dbg_mem_wdata,
	output         	o_dbg_mem_we,
	output         	o_dbg_data_access,
	output         	o_dbg_mem_read,
	output         	o_dbg_mem_write,
	output [31:0]   o_dbg_tmp
);

	parameter [0:0] BARREL_SHIFTER = 1;
	parameter [0:0] ENABLE_MULDIV = 1;
	parameter [0:0] ENABLE_COMPRESSED = 1;
	parameter [0:0] ENABLE_COUNTERS = 1;
	parameter [0:0] ENABLE_IRQ_QREGS = 0;

	parameter integer MEM_WORDS = 256;
	parameter [31:0] STACKADDR = 32'h 0000_0800;// (2*MEM_WORDS);       // end of memory
	parameter [31:0] PROGADDR_RESET = 32'h 0000_0000;
	parameter [31:0] PROGADDR_IRQ = 32'h 0020_0000;
	
	// picorv signals
	wire 		cpu_mem_valid;
	wire 		cpu_mem_instr;
	wire 		cpu_mem_ready;
	wire [31:0] cpu_mem_addr;
	wire [31:0] cpu_mem_wdata;
	wire [3:0] 	cpu_mem_wstrb;
	wire [31:0] cpu_mem_rdata;
	
	wire		cpu_read_request;
	wire		cpu_write_request;
	assign cpu_read_request = cpu_mem_instr || cpu_mem_wstrb == 4'b0;
	assign cpu_write_request = cpu_mem_wstrb != 4'b0;

// BEGIN DATA_DECL
reg [31 : 0] firmware[0 : 511];
reg [31 : 0] LanguageConstructsTestSource_SOC_Value;
reg [7 : 0] LanguageConstructsTestSource_SOC_Array[0 : 511];

// END DATA_DECL

// BEGIN DATA_CTRL
	// 32 bit memory logic for firmware
	wire 			firmware_ready;
	reg 			firmware_read_ready = 1'b0;
	reg 			firmware_write_ready = 1'b0;
	reg  [31:0] firmware_rdata = 32'b0;
	wire [31:0] firmware_wdata;	
	wire [31: 0]	firmware_address;
	wire 			firmware_we;
	reg  [1:0] 		firmware_write_state = 2'b0;
	wire 			firmware_address_valid;

	assign firmware_address_valid = cpu_mem_addr[31:20] == 12'h00;
	assign firmware_ready = firmware_read_ready || firmware_write_ready;
	
	assign firmware_wdata = {
		cpu_mem_wstrb[3] ? cpu_mem_wdata[31:24] : firmware_rdata[31:24],
		cpu_mem_wstrb[2] ? cpu_mem_wdata[23:16] : firmware_rdata[23:16],
		cpu_mem_wstrb[1] ? cpu_mem_wdata[15:8]  : firmware_rdata[15:8],
		cpu_mem_wstrb[0] ? cpu_mem_wdata[7:0]   : firmware_rdata[7:0]
	};

	assign firmware_we = firmware_write_state == 2'b1 && firmware_address_valid;
	assign firmware_address = cpu_mem_addr[31:2];
	
	always @(posedge clk)
	begin
		firmware_read_ready <= 1'b0;
		firmware_write_ready <= 1'b0;
		firmware_write_state <= 2'b0;
		firmware_rdata <= 32'b0;

		if (resetn && cpu_mem_valid && firmware_address_valid)
			begin	
				firmware_read_ready <= cpu_read_request;
				firmware_write_ready <= cpu_write_request && firmware_write_state == 2'b1;
			
				if (cpu_write_request)
				begin
					case (firmware_write_state)
						0: begin
							firmware_write_state <= 2'b1;
							// read ready in next cycle
						end
						1: begin
							firmware_write_state <= 2'b0;
						end
					endcase
				end
			end

		if (firmware_we)
			begin
				firmware[firmware_address] <= firmware_wdata;
			end

		firmware_rdata <= firmware[firmware_address];
	end

	wire 		LanguageConstructsTestSource_SOC_Value_ready;
	wire 		LanguageConstructsTestSource_SOC_Value_we;
	wire [31:0] LanguageConstructsTestSource_SOC_Value_wdata;	

	// byteenabled write
	assign LanguageConstructsTestSource_SOC_Value_wdata = {
		cpu_mem_wstrb[3] ? cpu_mem_wdata[31:24] : LanguageConstructsTestSource_SOC_Value[31:24],
		cpu_mem_wstrb[2] ? cpu_mem_wdata[23:16] : LanguageConstructsTestSource_SOC_Value[23:16],
		cpu_mem_wstrb[1] ? cpu_mem_wdata[15:8]  : LanguageConstructsTestSource_SOC_Value[15:8],
		cpu_mem_wstrb[0] ? cpu_mem_wdata[7:0]   : LanguageConstructsTestSource_SOC_Value[7:0]
	};
	
	assign LanguageConstructsTestSource_SOC_Value_ready = cpu_mem_addr[31:20] == 12'h800;
	assign LanguageConstructsTestSource_SOC_Value_we = LanguageConstructsTestSource_SOC_Value_ready && !cpu_mem_instr;
	
	// memory logic
	always @(posedge clk)
	begin
		if (resetn)
			begin
				if (LanguageConstructsTestSource_SOC_Value_we)
					begin
						LanguageConstructsTestSource_SOC_Value <= LanguageConstructsTestSource_SOC_Value_wdata;
					end
			end
		else
			begin
				LanguageConstructsTestSource_SOC_Value <= 32'b0;
			end
	end
	

	// 8 bit memory logic for LanguageConstructsTestSource_SOC_Array
	wire 			LanguageConstructsTestSource_SOC_Array_ready;
	reg 			LanguageConstructsTestSource_SOC_Array_read_ready = 0;
	reg 			LanguageConstructsTestSource_SOC_Array_write_ready = 0;
	reg  [31:0]		LanguageConstructsTestSource_SOC_Array_rdata = 0;
	reg  [7:0]		LanguageConstructsTestSource_SOC_Array_rdata_part = 0;
	wire [7:0]		LanguageConstructsTestSource_SOC_Array_wdata;	
	wire [31: 0]	LanguageConstructsTestSource_SOC_Array_read_address;
	wire [31: 0]	LanguageConstructsTestSource_SOC_Array_write_address;
	wire 			LanguageConstructsTestSource_SOC_Array_we;
	reg  [2:0] 		LanguageConstructsTestSource_SOC_Array_read_state = 0;
	wire 			LanguageConstructsTestSource_SOC_Array_address_valid;
	reg	 [1:0]		LanguageConstructsTestSource_SOC_Array_read_address_part = 0;
	wire [1:0]		LanguageConstructsTestSource_SOC_Array_write_address_part;

	assign o_dbg_tmp = LanguageConstructsTestSource_SOC_Array_rdata;

	assign LanguageConstructsTestSource_SOC_Array_address_valid = cpu_mem_addr[31:20] == 12'h801;
	assign LanguageConstructsTestSource_SOC_Array_ready = LanguageConstructsTestSource_SOC_Array_read_ready || LanguageConstructsTestSource_SOC_Array_write_ready;
	
	// could it be wrong? sure it can, but will deal later
	assign LanguageConstructsTestSource_SOC_Array_wdata = cpu_mem_wdata[7:0];

	assign LanguageConstructsTestSource_SOC_Array_we = cpu_write_request && cpu_mem_valid && LanguageConstructsTestSource_SOC_Array_address_valid;
	assign LanguageConstructsTestSource_SOC_Array_read_address = { cpu_mem_addr[31:2], LanguageConstructsTestSource_SOC_Array_read_address_part };
	assign LanguageConstructsTestSource_SOC_Array_write_address = { cpu_mem_addr[31:2], LanguageConstructsTestSource_SOC_Array_write_address_part };
	
	assign LanguageConstructsTestSource_SOC_Array_write_address_part = {
		cpu_mem_wstrb[3] ? 3 : 
		cpu_mem_wstrb[2] ? 2 :
		cpu_mem_wstrb[1] ? 1 :
		0 
	};

	always @(posedge clk)
	begin
		LanguageConstructsTestSource_SOC_Array_read_ready <= 1'b0;
		LanguageConstructsTestSource_SOC_Array_write_ready <= 1'b0;
		LanguageConstructsTestSource_SOC_Array_read_address_part <= 0;

		if (resetn && cpu_mem_valid && LanguageConstructsTestSource_SOC_Array_address_valid)
			begin	
				LanguageConstructsTestSource_SOC_Array_read_ready <= cpu_read_request && LanguageConstructsTestSource_SOC_Array_read_state == 3'b101;
				LanguageConstructsTestSource_SOC_Array_write_ready <= cpu_write_request;
			
				// 4 cycle read
				if (cpu_read_request && LanguageConstructsTestSource_SOC_Array_read_state <= 3'b101)
					begin
						LanguageConstructsTestSource_SOC_Array_read_state <= LanguageConstructsTestSource_SOC_Array_read_state + 1;
						if (LanguageConstructsTestSource_SOC_Array_read_state != 0)
							begin
								LanguageConstructsTestSource_SOC_Array_read_address_part <= LanguageConstructsTestSource_SOC_Array_read_address_part + 1;
								LanguageConstructsTestSource_SOC_Array_rdata <= { LanguageConstructsTestSource_SOC_Array_rdata_part, LanguageConstructsTestSource_SOC_Array_rdata[31:8] };
							end
					end
			end
		else
			begin
				LanguageConstructsTestSource_SOC_Array_read_state <= 0;
			end
	end

always @(posedge clk)
	begin
		LanguageConstructsTestSource_SOC_Array_rdata_part <= 0;

		if (resetn)
			begin
				if (LanguageConstructsTestSource_SOC_Array_we)
					begin
						LanguageConstructsTestSource_SOC_Array[LanguageConstructsTestSource_SOC_Array_write_address] <= LanguageConstructsTestSource_SOC_Array_wdata;
					end

				LanguageConstructsTestSource_SOC_Array_rdata_part <= LanguageConstructsTestSource_SOC_Array[LanguageConstructsTestSource_SOC_Array_read_address];
			end
	end

// END DATA_CTRL

	// feedback to cpu
	assign cpu_mem_ready = firmware_ready || LanguageConstructsTestSource_SOC_Value_ready || LanguageConstructsTestSource_SOC_Array_ready;
	assign cpu_mem_rdata = firmware_ready ? firmware_rdata : LanguageConstructsTestSource_SOC_Value_ready ? LanguageConstructsTestSource_SOC_Value : LanguageConstructsTestSource_SOC_Array_ready ? LanguageConstructsTestSource_SOC_Array_rdata : 32'b0;
		
	assign o_mem_valid = 	cpu_mem_valid;
	assign o_mem_instr = 	cpu_mem_instr;
	assign o_mem_addr = 	cpu_mem_addr;
	assign o_mem_wdata = 	cpu_mem_wdata;
	assign o_mem_wstrb = 	cpu_mem_wstrb;
	
	picorv32 #(
		.STACKADDR(STACKADDR),
		.PROGADDR_RESET(PROGADDR_RESET),
		.PROGADDR_IRQ(PROGADDR_IRQ),
		.BARREL_SHIFTER(BARREL_SHIFTER),
		.COMPRESSED_ISA(ENABLE_COMPRESSED),
		.ENABLE_COUNTERS(ENABLE_COUNTERS),
		.ENABLE_MUL(ENABLE_MULDIV),
		.ENABLE_DIV(ENABLE_MULDIV),
		.ENABLE_IRQ(1),
		.ENABLE_IRQ_QREGS(ENABLE_IRQ_QREGS)
	) cpu (
		.clk         (clk        	),
		.resetn      (resetn     	),
		.mem_valid   (cpu_mem_valid ),
		.mem_instr   (cpu_mem_instr ),
		.mem_ready   (cpu_mem_ready ),
		.mem_addr    (cpu_mem_addr  ),
		.mem_wdata   (cpu_mem_wdata ),
		.mem_wstrb   (cpu_mem_wstrb ),
		.mem_rdata   (cpu_mem_rdata ),
		.irq         (0        	 	)
	);
	
	// connect debug and diagnostics
			
	assign o_dbg_mem_valid = firmware_ready;
	assign o_dbg_mem_rdata = firmware_rdata;
	assign o_dbg_mem_wdata = firmware_wdata;
	assign o_dbg_mem_we = firmware_we;

	//assign o_dbg_mem_rdata = data_rdata_part;
	//assign o_dbg_mem_wdata = data_read_address_part;
	//assign o_dbg_mem_we = data_we;
	
	//assign o_dbg_data_access = data_address_valid;
	assign o_dbg_mem_read = cpu_read_request;
	assign o_dbg_mem_write = cpu_write_request;
	
	initial
	begin
// BEGIN MEM_INIT
/*000*/firmware[0] = 32'h1740006F;
/*004*/firmware[1] = 32'h00000013;
/*008*/firmware[2] = 32'h00000013;
/*00C*/firmware[3] = 32'h00000013;
/*010*/firmware[4] = 32'h00102223;
/*014*/firmware[5] = 32'h00202423;
/*018*/firmware[6] = 32'h0000408B;
/*01C*/firmware[7] = 32'h00102623;
/*020*/firmware[8] = 32'h0000C08B;
/*024*/firmware[9] = 32'h00102823;
/*028*/firmware[10] = 32'h00001137;
/*02C*/firmware[11] = 32'hF8010113;
/*030*/firmware[12] = 32'h0000408B;
/*034*/firmware[13] = 32'h00112023;
/*038*/firmware[14] = 32'h00402083;
/*03C*/firmware[15] = 32'h00112223;
/*040*/firmware[16] = 32'h00802083;
/*044*/firmware[17] = 32'h00112423;
/*048*/firmware[18] = 32'h00312623;
/*04C*/firmware[19] = 32'h00412823;
/*050*/firmware[20] = 32'h00512A23;
/*054*/firmware[21] = 32'h00612C23;
/*058*/firmware[22] = 32'h00712E23;
/*05C*/firmware[23] = 32'h02812023;
/*060*/firmware[24] = 32'h02912223;
/*064*/firmware[25] = 32'h02A12423;
/*068*/firmware[26] = 32'h02B12623;
/*06C*/firmware[27] = 32'h02C12823;
/*070*/firmware[28] = 32'h02D12A23;
/*074*/firmware[29] = 32'h02E12C23;
/*078*/firmware[30] = 32'h02F12E23;
/*07C*/firmware[31] = 32'h05012023;
/*080*/firmware[32] = 32'h05112223;
/*084*/firmware[33] = 32'h05212423;
/*088*/firmware[34] = 32'h05312623;
/*08C*/firmware[35] = 32'h05412823;
/*090*/firmware[36] = 32'h05512A23;
/*094*/firmware[37] = 32'h05612C23;
/*098*/firmware[38] = 32'h05712E23;
/*09C*/firmware[39] = 32'h07812023;
/*0A0*/firmware[40] = 32'h07912223;
/*0A4*/firmware[41] = 32'h07A12423;
/*0A8*/firmware[42] = 32'h07B12623;
/*0AC*/firmware[43] = 32'h07C12823;
/*0B0*/firmware[44] = 32'h07D12A23;
/*0B4*/firmware[45] = 32'h07E12C23;
/*0B8*/firmware[46] = 32'h07F12E23;
/*0BC*/firmware[47] = 32'h0000C50B;
/*0C0*/firmware[48] = 32'h00010593;
/*0C4*/firmware[49] = 32'h00002083;
/*0C8*/firmware[50] = 32'h00100463;
/*0CC*/firmware[51] = 32'h000080E7;
/*0D0*/firmware[52] = 32'h00012083;
/*0D4*/firmware[53] = 32'h0200A00B;
/*0D8*/firmware[54] = 32'h00412083;
/*0DC*/firmware[55] = 32'h0200A08B;
/*0E0*/firmware[56] = 32'h00812083;
/*0E4*/firmware[57] = 32'h00102223;
/*0E8*/firmware[58] = 32'h00C12183;
/*0EC*/firmware[59] = 32'h01012203;
/*0F0*/firmware[60] = 32'h01412283;
/*0F4*/firmware[61] = 32'h01812303;
/*0F8*/firmware[62] = 32'h01C12383;
/*0FC*/firmware[63] = 32'h02012403;
/*100*/firmware[64] = 32'h02412483;
/*104*/firmware[65] = 32'h02812503;
/*108*/firmware[66] = 32'h02C12583;
/*10C*/firmware[67] = 32'h03012603;
/*110*/firmware[68] = 32'h03412683;
/*114*/firmware[69] = 32'h03812703;
/*118*/firmware[70] = 32'h03C12783;
/*11C*/firmware[71] = 32'h04012803;
/*120*/firmware[72] = 32'h04412883;
/*124*/firmware[73] = 32'h04812903;
/*128*/firmware[74] = 32'h04C12983;
/*12C*/firmware[75] = 32'h05012A03;
/*130*/firmware[76] = 32'h05412A83;
/*134*/firmware[77] = 32'h05812B03;
/*138*/firmware[78] = 32'h05C12B83;
/*13C*/firmware[79] = 32'h06012C03;
/*140*/firmware[80] = 32'h06412C83;
/*144*/firmware[81] = 32'h06812D03;
/*148*/firmware[82] = 32'h06C12D83;
/*14C*/firmware[83] = 32'h07012E03;
/*150*/firmware[84] = 32'h07412E83;
/*154*/firmware[85] = 32'h07812F03;
/*158*/firmware[86] = 32'h07C12F83;
/*15C*/firmware[87] = 32'h0000C08B;
/*160*/firmware[88] = 32'h00402103;
/*164*/firmware[89] = 32'h00000013;
/*168*/firmware[90] = 32'h00000013;
/*16C*/firmware[91] = 32'h00000013;
/*170*/firmware[92] = 32'h0400000B;
/*174*/firmware[93] = 32'h00000093;
/*178*/firmware[94] = 32'h00000193;
/*17C*/firmware[95] = 32'h00000213;
/*180*/firmware[96] = 32'h00000293;
/*184*/firmware[97] = 32'h00000313;
/*188*/firmware[98] = 32'h00000393;
/*18C*/firmware[99] = 32'h00000413;
/*190*/firmware[100] = 32'h00000493;
/*194*/firmware[101] = 32'h00000513;
/*198*/firmware[102] = 32'h00000593;
/*19C*/firmware[103] = 32'h00000613;
/*1A0*/firmware[104] = 32'h00000693;
/*1A4*/firmware[105] = 32'h00000713;
/*1A8*/firmware[106] = 32'h00000793;
/*1AC*/firmware[107] = 32'h00000813;
/*1B0*/firmware[108] = 32'h00000893;
/*1B4*/firmware[109] = 32'h00000913;
/*1B8*/firmware[110] = 32'h00000993;
/*1BC*/firmware[111] = 32'h00000A13;
/*1C0*/firmware[112] = 32'h00000A93;
/*1C4*/firmware[113] = 32'h00000B13;
/*1C8*/firmware[114] = 32'h00000B93;
/*1CC*/firmware[115] = 32'h00000C13;
/*1D0*/firmware[116] = 32'h00000C93;
/*1D4*/firmware[117] = 32'h00000D13;
/*1D8*/firmware[118] = 32'h00000D93;
/*1DC*/firmware[119] = 32'h00000E13;
/*1E0*/firmware[120] = 32'h00000E93;
/*1E4*/firmware[121] = 32'h00000F13;
/*1E8*/firmware[122] = 32'h00000F93;
/*1EC*/firmware[123] = 32'h018000EF;
/*1F0*/firmware[124] = 32'h0000006F;
/*1F4*/firmware[125] = 32'h00000000;
/*1F8*/firmware[126] = 32'h00000000;
/*1FC*/firmware[127] = 32'h0605650B;
/*200*/firmware[128] = 32'h00008067;
/*204*/firmware[129] = 32'hFE010113;
/*208*/firmware[130] = 32'h00112E23;
/*20C*/firmware[131] = 32'h00812C23;
/*210*/firmware[132] = 32'h02010413;
/*214*/firmware[133] = 32'h0FF00513;
/*218*/firmware[134] = 32'hFE5FF0EF;
/*21C*/firmware[135] = 32'h59C00793;
/*220*/firmware[136] = 32'hFEF42623;
/*224*/firmware[137] = 32'hFEC42703;
/*228*/firmware[138] = 32'h59C00793;
/*22C*/firmware[139] = 32'h00F77C63;
/*230*/firmware[140] = 32'hFEC42783;
/*234*/firmware[141] = 32'h00478713;
/*238*/firmware[142] = 32'hFEE42623;
/*23C*/firmware[143] = 32'h0007A023;
/*240*/firmware[144] = 32'hFE5FF06F;
/*244*/firmware[145] = 32'h210000EF;
/*248*/firmware[146] = 32'h00000013;
/*24C*/firmware[147] = 32'h01C12083;
/*250*/firmware[148] = 32'h01812403;
/*254*/firmware[149] = 32'h02010113;
/*258*/firmware[150] = 32'h00008067;
/*25C*/firmware[151] = 32'hFE010113;
/*260*/firmware[152] = 32'h00812E23;
/*264*/firmware[153] = 32'h02010413;
/*268*/firmware[154] = 32'hFEA42623;
/*26C*/firmware[155] = 32'hFEC42703;
/*270*/firmware[156] = 32'h00400793;
/*274*/firmware[157] = 32'h00E7C863;
/*278*/firmware[158] = 32'h800007B7;
/*27C*/firmware[159] = 32'h0007A023;
/*280*/firmware[160] = 32'h0300006F;
/*284*/firmware[161] = 32'hFEC42703;
/*288*/firmware[162] = 32'h00700793;
/*28C*/firmware[163] = 32'h00E7CA63;
/*290*/firmware[164] = 32'h800007B7;
/*294*/firmware[165] = 32'h00100713;
/*298*/firmware[166] = 32'h00E7A023;
/*29C*/firmware[167] = 32'h0140006F;
/*2A0*/firmware[168] = 32'h800007B7;
/*2A4*/firmware[169] = 32'hFEC42703;
/*2A8*/firmware[170] = 32'h00A70713;
/*2AC*/firmware[171] = 32'h00E7A023;
/*2B0*/firmware[172] = 32'h00000013;
/*2B4*/firmware[173] = 32'h01C12403;
/*2B8*/firmware[174] = 32'h02010113;
/*2BC*/firmware[175] = 32'h00008067;
/*2C0*/firmware[176] = 32'hFE010113;
/*2C4*/firmware[177] = 32'h00812E23;
/*2C8*/firmware[178] = 32'h02010413;
/*2CC*/firmware[179] = 32'hFEA42623;
/*2D0*/firmware[180] = 32'hFEC42703;
/*2D4*/firmware[181] = 32'h00100793;
/*2D8*/firmware[182] = 32'h02F70C63;
/*2DC*/firmware[183] = 32'hFEC42703;
/*2E0*/firmware[184] = 32'h00100793;
/*2E4*/firmware[185] = 32'h00E7C863;
/*2E8*/firmware[186] = 32'hFEC42783;
/*2EC*/firmware[187] = 32'h00078C63;
/*2F0*/firmware[188] = 32'h03C0006F;
/*2F4*/firmware[189] = 32'hFEC42703;
/*2F8*/firmware[190] = 32'h00300793;
/*2FC*/firmware[191] = 32'h02E7C863;
/*300*/firmware[192] = 32'h01C0006F;
/*304*/firmware[193] = 32'h800007B7;
/*308*/firmware[194] = 32'h0007A023;
/*30C*/firmware[195] = 32'h03C0006F;
/*310*/firmware[196] = 32'h800007B7;
/*314*/firmware[197] = 32'h0007A023;
/*318*/firmware[198] = 32'h0300006F;
/*31C*/firmware[199] = 32'h800007B7;
/*320*/firmware[200] = 32'h00200713;
/*324*/firmware[201] = 32'h00E7A023;
/*328*/firmware[202] = 32'h0200006F;
/*32C*/firmware[203] = 32'h800006B7;
/*330*/firmware[204] = 32'hFEC42703;
/*334*/firmware[205] = 32'h00070793;
/*338*/firmware[206] = 32'h00179793;
/*33C*/firmware[207] = 32'h00E787B3;
/*340*/firmware[208] = 32'h00F6A023;
/*344*/firmware[209] = 32'h00000013;
/*348*/firmware[210] = 32'h00000013;
/*34C*/firmware[211] = 32'h01C12403;
/*350*/firmware[212] = 32'h02010113;
/*354*/firmware[213] = 32'h00008067;
/*358*/firmware[214] = 32'hFD010113;
/*35C*/firmware[215] = 32'h02812623;
/*360*/firmware[216] = 32'h03010413;
/*364*/firmware[217] = 32'hFCA42E23;
/*368*/firmware[218] = 32'hFE042623;
/*36C*/firmware[219] = 32'hFEC42703;
/*370*/firmware[220] = 32'hFDC42783;
/*374*/firmware[221] = 32'h02F75663;
/*378*/firmware[222] = 32'h800007B7;
/*37C*/firmware[223] = 32'h0007A683;
/*380*/firmware[224] = 32'h800007B7;
/*384*/firmware[225] = 32'hFEC42703;
/*388*/firmware[226] = 32'h02E68733;
/*38C*/firmware[227] = 32'h00E7A023;
/*390*/firmware[228] = 32'hFEC42783;
/*394*/firmware[229] = 32'h00178793;
/*398*/firmware[230] = 32'hFEF42623;
/*39C*/firmware[231] = 32'hFD1FF06F;
/*3A0*/firmware[232] = 32'hFDC42783;
/*3A4*/firmware[233] = 32'hFEF42423;
/*3A8*/firmware[234] = 32'hFE842783;
/*3AC*/firmware[235] = 32'h0207C663;
/*3B0*/firmware[236] = 32'h800007B7;
/*3B4*/firmware[237] = 32'h0007A683;
/*3B8*/firmware[238] = 32'h800007B7;
/*3BC*/firmware[239] = 32'hFE842703;
/*3C0*/firmware[240] = 32'h02E6C733;
/*3C4*/firmware[241] = 32'h00E7A023;
/*3C8*/firmware[242] = 32'hFE842783;
/*3CC*/firmware[243] = 32'hFFF78793;
/*3D0*/firmware[244] = 32'hFEF42423;
/*3D4*/firmware[245] = 32'hFD5FF06F;
/*3D8*/firmware[246] = 32'hFDC42783;
/*3DC*/firmware[247] = 32'hFFF78713;
/*3E0*/firmware[248] = 32'hFCE42E23;
/*3E4*/firmware[249] = 32'hFFF7C793;
/*3E8*/firmware[250] = 32'h01F7D793;
/*3EC*/firmware[251] = 32'h0FF7F793;
/*3F0*/firmware[252] = 32'h02078063;
/*3F4*/firmware[253] = 32'h800007B7;
/*3F8*/firmware[254] = 32'h0007A683;
/*3FC*/firmware[255] = 32'h800007B7;
/*400*/firmware[256] = 32'hFDC42703;
/*404*/firmware[257] = 32'h00E68733;
/*408*/firmware[258] = 32'h00E7A023;
/*40C*/firmware[259] = 32'hFCDFF06F;
/*410*/firmware[260] = 32'h800007B7;
/*414*/firmware[261] = 32'h0007A683;
/*418*/firmware[262] = 32'h800007B7;
/*41C*/firmware[263] = 32'hFDC42703;
/*420*/firmware[264] = 32'h00E68733;
/*424*/firmware[265] = 32'h00E7A023;
/*428*/firmware[266] = 32'hFDC42783;
/*42C*/firmware[267] = 32'h00178713;
/*430*/firmware[268] = 32'hFCE42E23;
/*434*/firmware[269] = 32'h00A7A793;
/*438*/firmware[270] = 32'h0FF7F793;
/*43C*/firmware[271] = 32'h00078463;
/*440*/firmware[272] = 32'hFD1FF06F;
/*444*/firmware[273] = 32'h00000013;
/*448*/firmware[274] = 32'h02C12403;
/*44C*/firmware[275] = 32'h03010113;
/*450*/firmware[276] = 32'h00008067;
/*454*/firmware[277] = 32'hFE010113;
/*458*/firmware[278] = 32'h00112E23;
/*45C*/firmware[279] = 32'h00812C23;
/*460*/firmware[280] = 32'h02010413;
/*464*/firmware[281] = 32'hFE042623;
/*468*/firmware[282] = 32'hFEC42703;
/*46C*/firmware[283] = 32'h00900793;
/*470*/firmware[284] = 32'h02E7C063;
/*474*/firmware[285] = 32'hFEC42503;
/*478*/firmware[286] = 32'hDE5FF0EF;
/*47C*/firmware[287] = 32'hFEC42503;
/*480*/firmware[288] = 32'hE41FF0EF;
/*484*/firmware[289] = 32'hFEC42503;
/*488*/firmware[290] = 32'hED1FF0EF;
/*48C*/firmware[291] = 32'hFDDFF06F;
/*490*/firmware[292] = 32'h00000013;
/*494*/firmware[293] = 32'h01C12083;
/*498*/firmware[294] = 32'h01812403;
/*49C*/firmware[295] = 32'h02010113;
/*4A0*/firmware[296] = 32'h00008067;
/*4A4*/firmware[297] = 32'h00000010;
/*4A8*/firmware[298] = 32'h00000000;
/*4AC*/firmware[299] = 32'h00527A01;
/*4B0*/firmware[300] = 32'h01017C01;
/*4B4*/firmware[301] = 32'h00020D1B;
/*4B8*/firmware[302] = 32'h00000024;
/*4BC*/firmware[303] = 32'h00000018;
/*4C0*/firmware[304] = 32'hFFFFFD44;
/*4C4*/firmware[305] = 32'h00000058;
/*4C8*/firmware[306] = 32'h200E4400;
/*4CC*/firmware[307] = 32'h88018148;
/*4D0*/firmware[308] = 32'h080C4402;
/*4D4*/firmware[309] = 32'hC13C0200;
/*4D8*/firmware[310] = 32'h0D44C844;
/*4DC*/firmware[311] = 32'h00000002;
/*4E0*/firmware[312] = 32'h00000010;
/*4E4*/firmware[313] = 32'h00000000;
/*4E8*/firmware[314] = 32'h00527A01;
/*4EC*/firmware[315] = 32'h01017C01;
/*4F0*/firmware[316] = 32'h00020D1B;
/*4F4*/firmware[317] = 32'h00000020;
/*4F8*/firmware[318] = 32'h00000018;
/*4FC*/firmware[319] = 32'hFFFFFD60;
/*500*/firmware[320] = 32'h00000064;
/*504*/firmware[321] = 32'h200E4400;
/*508*/firmware[322] = 32'h44018844;
/*50C*/firmware[323] = 32'h0200080C;
/*510*/firmware[324] = 32'h0D44C850;
/*514*/firmware[325] = 32'h00000002;
/*518*/firmware[326] = 32'h00000020;
/*51C*/firmware[327] = 32'h0000003C;
/*520*/firmware[328] = 32'hFFFFFDA0;
/*524*/firmware[329] = 32'h00000098;
/*528*/firmware[330] = 32'h200E4400;
/*52C*/firmware[331] = 32'h44018844;
/*530*/firmware[332] = 32'h0200080C;
/*534*/firmware[333] = 32'h0D44C884;
/*538*/firmware[334] = 32'h00000002;
/*53C*/firmware[335] = 32'h00000020;
/*540*/firmware[336] = 32'h00000060;
/*544*/firmware[337] = 32'hFFFFFE14;
/*548*/firmware[338] = 32'h000000FC;
/*54C*/firmware[339] = 32'h300E4400;
/*550*/firmware[340] = 32'h44018844;
/*554*/firmware[341] = 32'h0200080C;
/*558*/firmware[342] = 32'h0D44C8E8;
/*55C*/firmware[343] = 32'h00000002;
/*560*/firmware[344] = 32'h00000024;
/*564*/firmware[345] = 32'h00000084;
/*568*/firmware[346] = 32'hFFFFFEEC;
/*56C*/firmware[347] = 32'h00000050;
/*570*/firmware[348] = 32'h200E4400;
/*574*/firmware[349] = 32'h88018148;
/*578*/firmware[350] = 32'h080C4402;
/*57C*/firmware[351] = 32'hC1340200;
/*580*/firmware[352] = 32'h0D44C844;
/*584*/firmware[353] = 32'h00000002;
/*588*/firmware[354] = 32'h00000000;
/*58C*/firmware[355] = 32'h00000000;
/*590*/firmware[356] = 32'h00000000;
/*594*/firmware[357] = 32'h00000000;
/*598*/firmware[358] = 32'h00000000;
/*59C*/firmware[359] = 32'h00000000;
/*5A0*/firmware[360] = 32'h00000000;
/*5A4*/firmware[361] = 32'h00000000;
/*5A8*/firmware[362] = 32'h00000000;
/*5AC*/firmware[363] = 32'h00000000;
/*5B0*/firmware[364] = 32'h00000000;
/*5B4*/firmware[365] = 32'h00000000;
/*5B8*/firmware[366] = 32'h00000000;
/*5BC*/firmware[367] = 32'h00000000;
/*5C0*/firmware[368] = 32'h00000000;
/*5C4*/firmware[369] = 32'h00000000;
/*5C8*/firmware[370] = 32'h00000000;
/*5CC*/firmware[371] = 32'h00000000;
/*5D0*/firmware[372] = 32'h00000000;
/*5D4*/firmware[373] = 32'h00000000;
/*5D8*/firmware[374] = 32'h00000000;
/*5DC*/firmware[375] = 32'h00000000;
/*5E0*/firmware[376] = 32'h00000000;
/*5E4*/firmware[377] = 32'h00000000;
/*5E8*/firmware[378] = 32'h00000000;
/*5EC*/firmware[379] = 32'h00000000;
/*5F0*/firmware[380] = 32'h00000000;
/*5F4*/firmware[381] = 32'h00000000;
/*5F8*/firmware[382] = 32'h00000000;
/*5FC*/firmware[383] = 32'h00000000;
/*600*/firmware[384] = 32'h00000000;
/*604*/firmware[385] = 32'h00000000;
/*608*/firmware[386] = 32'h00000000;
/*60C*/firmware[387] = 32'h00000000;
/*610*/firmware[388] = 32'h00000000;
/*614*/firmware[389] = 32'h00000000;
/*618*/firmware[390] = 32'h00000000;
/*61C*/firmware[391] = 32'h00000000;
/*620*/firmware[392] = 32'h00000000;
/*624*/firmware[393] = 32'h00000000;
/*628*/firmware[394] = 32'h00000000;
/*62C*/firmware[395] = 32'h00000000;
/*630*/firmware[396] = 32'h00000000;
/*634*/firmware[397] = 32'h00000000;
/*638*/firmware[398] = 32'h00000000;
/*63C*/firmware[399] = 32'h00000000;
/*640*/firmware[400] = 32'h00000000;
/*644*/firmware[401] = 32'h00000000;
/*648*/firmware[402] = 32'h00000000;
/*64C*/firmware[403] = 32'h00000000;
/*650*/firmware[404] = 32'h00000000;
/*654*/firmware[405] = 32'h00000000;
/*658*/firmware[406] = 32'h00000000;
/*65C*/firmware[407] = 32'h00000000;
/*660*/firmware[408] = 32'h00000000;
/*664*/firmware[409] = 32'h00000000;
/*668*/firmware[410] = 32'h00000000;
/*66C*/firmware[411] = 32'h00000000;
/*670*/firmware[412] = 32'h00000000;
/*674*/firmware[413] = 32'h00000000;
/*678*/firmware[414] = 32'h00000000;
/*67C*/firmware[415] = 32'h00000000;
/*680*/firmware[416] = 32'h00000000;
/*684*/firmware[417] = 32'h00000000;
/*688*/firmware[418] = 32'h00000000;
/*68C*/firmware[419] = 32'h00000000;
/*690*/firmware[420] = 32'h00000000;
/*694*/firmware[421] = 32'h00000000;
/*698*/firmware[422] = 32'h00000000;
/*69C*/firmware[423] = 32'h00000000;
/*6A0*/firmware[424] = 32'h00000000;
/*6A4*/firmware[425] = 32'h00000000;
/*6A8*/firmware[426] = 32'h00000000;
/*6AC*/firmware[427] = 32'h00000000;
/*6B0*/firmware[428] = 32'h00000000;
/*6B4*/firmware[429] = 32'h00000000;
/*6B8*/firmware[430] = 32'h00000000;
/*6BC*/firmware[431] = 32'h00000000;
/*6C0*/firmware[432] = 32'h00000000;
/*6C4*/firmware[433] = 32'h00000000;
/*6C8*/firmware[434] = 32'h00000000;
/*6CC*/firmware[435] = 32'h00000000;
/*6D0*/firmware[436] = 32'h00000000;
/*6D4*/firmware[437] = 32'h00000000;
/*6D8*/firmware[438] = 32'h00000000;
/*6DC*/firmware[439] = 32'h00000000;
/*6E0*/firmware[440] = 32'h00000000;
/*6E4*/firmware[441] = 32'h00000000;
/*6E8*/firmware[442] = 32'h00000000;
/*6EC*/firmware[443] = 32'h00000000;
/*6F0*/firmware[444] = 32'h00000000;
/*6F4*/firmware[445] = 32'h00000000;
/*6F8*/firmware[446] = 32'h00000000;
/*6FC*/firmware[447] = 32'h00000000;
/*700*/firmware[448] = 32'h00000000;
/*704*/firmware[449] = 32'h00000000;
/*708*/firmware[450] = 32'h00000000;
/*70C*/firmware[451] = 32'h00000000;
/*710*/firmware[452] = 32'h00000000;
/*714*/firmware[453] = 32'h00000000;
/*718*/firmware[454] = 32'h00000000;
/*71C*/firmware[455] = 32'h00000000;
/*720*/firmware[456] = 32'h00000000;
/*724*/firmware[457] = 32'h00000000;
/*728*/firmware[458] = 32'h00000000;
/*72C*/firmware[459] = 32'h00000000;
/*730*/firmware[460] = 32'h00000000;
/*734*/firmware[461] = 32'h00000000;
/*738*/firmware[462] = 32'h00000000;
/*73C*/firmware[463] = 32'h00000000;
/*740*/firmware[464] = 32'h00000000;
/*744*/firmware[465] = 32'h00000000;
/*748*/firmware[466] = 32'h00000000;
/*74C*/firmware[467] = 32'h00000000;
/*750*/firmware[468] = 32'h00000000;
/*754*/firmware[469] = 32'h00000000;
/*758*/firmware[470] = 32'h00000000;
/*75C*/firmware[471] = 32'h00000000;
/*760*/firmware[472] = 32'h00000000;
/*764*/firmware[473] = 32'h00000000;
/*768*/firmware[474] = 32'h00000000;
/*76C*/firmware[475] = 32'h00000000;
/*770*/firmware[476] = 32'h00000000;
/*774*/firmware[477] = 32'h00000000;
/*778*/firmware[478] = 32'h00000000;
/*77C*/firmware[479] = 32'h00000000;
/*780*/firmware[480] = 32'h00000000;
/*784*/firmware[481] = 32'h00000000;
/*788*/firmware[482] = 32'h00000000;
/*78C*/firmware[483] = 32'h00000000;
/*790*/firmware[484] = 32'h00000000;
/*794*/firmware[485] = 32'h00000000;
/*798*/firmware[486] = 32'h00000000;
/*79C*/firmware[487] = 32'h00000000;
/*7A0*/firmware[488] = 32'h00000000;
/*7A4*/firmware[489] = 32'h00000000;
/*7A8*/firmware[490] = 32'h00000000;
/*7AC*/firmware[491] = 32'h00000000;
/*7B0*/firmware[492] = 32'h00000000;
/*7B4*/firmware[493] = 32'h00000000;
/*7B8*/firmware[494] = 32'h00000000;
/*7BC*/firmware[495] = 32'h00000000;
/*7C0*/firmware[496] = 32'h00000000;
/*7C4*/firmware[497] = 32'h00000000;
/*7C8*/firmware[498] = 32'h00000000;
/*7CC*/firmware[499] = 32'h00000000;
/*7D0*/firmware[500] = 32'h00000000;
/*7D4*/firmware[501] = 32'h00000000;
/*7D8*/firmware[502] = 32'h00000000;
/*7DC*/firmware[503] = 32'h00000000;
/*7E0*/firmware[504] = 32'h00000000;
/*7E4*/firmware[505] = 32'h00000000;
/*7E8*/firmware[506] = 32'h00000000;
/*7EC*/firmware[507] = 32'h00000000;
/*7F0*/firmware[508] = 32'h00000000;
/*7F4*/firmware[509] = 32'h00000000;
/*7F8*/firmware[510] = 32'h00000000;
/*7FC*/firmware[511] = 32'h00000000;
/*000*/LanguageConstructsTestSource_SOC_Array[0] = 8'h00;
/*001*/LanguageConstructsTestSource_SOC_Array[1] = 8'h00;
/*002*/LanguageConstructsTestSource_SOC_Array[2] = 8'h00;
/*003*/LanguageConstructsTestSource_SOC_Array[3] = 8'h00;
/*004*/LanguageConstructsTestSource_SOC_Array[4] = 8'h00;
/*005*/LanguageConstructsTestSource_SOC_Array[5] = 8'h00;
/*006*/LanguageConstructsTestSource_SOC_Array[6] = 8'h00;
/*007*/LanguageConstructsTestSource_SOC_Array[7] = 8'h00;
/*008*/LanguageConstructsTestSource_SOC_Array[8] = 8'h00;
/*009*/LanguageConstructsTestSource_SOC_Array[9] = 8'h00;
/*00A*/LanguageConstructsTestSource_SOC_Array[10] = 8'h00;
/*00B*/LanguageConstructsTestSource_SOC_Array[11] = 8'h00;
/*00C*/LanguageConstructsTestSource_SOC_Array[12] = 8'h00;
/*00D*/LanguageConstructsTestSource_SOC_Array[13] = 8'h00;
/*00E*/LanguageConstructsTestSource_SOC_Array[14] = 8'h00;
/*00F*/LanguageConstructsTestSource_SOC_Array[15] = 8'h00;
/*010*/LanguageConstructsTestSource_SOC_Array[16] = 8'h00;
/*011*/LanguageConstructsTestSource_SOC_Array[17] = 8'h00;
/*012*/LanguageConstructsTestSource_SOC_Array[18] = 8'h00;
/*013*/LanguageConstructsTestSource_SOC_Array[19] = 8'h00;
/*014*/LanguageConstructsTestSource_SOC_Array[20] = 8'h00;
/*015*/LanguageConstructsTestSource_SOC_Array[21] = 8'h00;
/*016*/LanguageConstructsTestSource_SOC_Array[22] = 8'h00;
/*017*/LanguageConstructsTestSource_SOC_Array[23] = 8'h00;
/*018*/LanguageConstructsTestSource_SOC_Array[24] = 8'h00;
/*019*/LanguageConstructsTestSource_SOC_Array[25] = 8'h00;
/*01A*/LanguageConstructsTestSource_SOC_Array[26] = 8'h00;
/*01B*/LanguageConstructsTestSource_SOC_Array[27] = 8'h00;
/*01C*/LanguageConstructsTestSource_SOC_Array[28] = 8'h00;
/*01D*/LanguageConstructsTestSource_SOC_Array[29] = 8'h00;
/*01E*/LanguageConstructsTestSource_SOC_Array[30] = 8'h00;
/*01F*/LanguageConstructsTestSource_SOC_Array[31] = 8'h00;
/*020*/LanguageConstructsTestSource_SOC_Array[32] = 8'h00;
/*021*/LanguageConstructsTestSource_SOC_Array[33] = 8'h00;
/*022*/LanguageConstructsTestSource_SOC_Array[34] = 8'h00;
/*023*/LanguageConstructsTestSource_SOC_Array[35] = 8'h00;
/*024*/LanguageConstructsTestSource_SOC_Array[36] = 8'h00;
/*025*/LanguageConstructsTestSource_SOC_Array[37] = 8'h00;
/*026*/LanguageConstructsTestSource_SOC_Array[38] = 8'h00;
/*027*/LanguageConstructsTestSource_SOC_Array[39] = 8'h00;
/*028*/LanguageConstructsTestSource_SOC_Array[40] = 8'h00;
/*029*/LanguageConstructsTestSource_SOC_Array[41] = 8'h00;
/*02A*/LanguageConstructsTestSource_SOC_Array[42] = 8'h00;
/*02B*/LanguageConstructsTestSource_SOC_Array[43] = 8'h00;
/*02C*/LanguageConstructsTestSource_SOC_Array[44] = 8'h00;
/*02D*/LanguageConstructsTestSource_SOC_Array[45] = 8'h00;
/*02E*/LanguageConstructsTestSource_SOC_Array[46] = 8'h00;
/*02F*/LanguageConstructsTestSource_SOC_Array[47] = 8'h00;
/*030*/LanguageConstructsTestSource_SOC_Array[48] = 8'h00;
/*031*/LanguageConstructsTestSource_SOC_Array[49] = 8'h00;
/*032*/LanguageConstructsTestSource_SOC_Array[50] = 8'h00;
/*033*/LanguageConstructsTestSource_SOC_Array[51] = 8'h00;
/*034*/LanguageConstructsTestSource_SOC_Array[52] = 8'h00;
/*035*/LanguageConstructsTestSource_SOC_Array[53] = 8'h00;
/*036*/LanguageConstructsTestSource_SOC_Array[54] = 8'h00;
/*037*/LanguageConstructsTestSource_SOC_Array[55] = 8'h00;
/*038*/LanguageConstructsTestSource_SOC_Array[56] = 8'h00;
/*039*/LanguageConstructsTestSource_SOC_Array[57] = 8'h00;
/*03A*/LanguageConstructsTestSource_SOC_Array[58] = 8'h00;
/*03B*/LanguageConstructsTestSource_SOC_Array[59] = 8'h00;
/*03C*/LanguageConstructsTestSource_SOC_Array[60] = 8'h00;
/*03D*/LanguageConstructsTestSource_SOC_Array[61] = 8'h00;
/*03E*/LanguageConstructsTestSource_SOC_Array[62] = 8'h00;
/*03F*/LanguageConstructsTestSource_SOC_Array[63] = 8'h00;
/*040*/LanguageConstructsTestSource_SOC_Array[64] = 8'h00;
/*041*/LanguageConstructsTestSource_SOC_Array[65] = 8'h00;
/*042*/LanguageConstructsTestSource_SOC_Array[66] = 8'h00;
/*043*/LanguageConstructsTestSource_SOC_Array[67] = 8'h00;
/*044*/LanguageConstructsTestSource_SOC_Array[68] = 8'h00;
/*045*/LanguageConstructsTestSource_SOC_Array[69] = 8'h00;
/*046*/LanguageConstructsTestSource_SOC_Array[70] = 8'h00;
/*047*/LanguageConstructsTestSource_SOC_Array[71] = 8'h00;
/*048*/LanguageConstructsTestSource_SOC_Array[72] = 8'h00;
/*049*/LanguageConstructsTestSource_SOC_Array[73] = 8'h00;
/*04A*/LanguageConstructsTestSource_SOC_Array[74] = 8'h00;
/*04B*/LanguageConstructsTestSource_SOC_Array[75] = 8'h00;
/*04C*/LanguageConstructsTestSource_SOC_Array[76] = 8'h00;
/*04D*/LanguageConstructsTestSource_SOC_Array[77] = 8'h00;
/*04E*/LanguageConstructsTestSource_SOC_Array[78] = 8'h00;
/*04F*/LanguageConstructsTestSource_SOC_Array[79] = 8'h00;
/*050*/LanguageConstructsTestSource_SOC_Array[80] = 8'h00;
/*051*/LanguageConstructsTestSource_SOC_Array[81] = 8'h00;
/*052*/LanguageConstructsTestSource_SOC_Array[82] = 8'h00;
/*053*/LanguageConstructsTestSource_SOC_Array[83] = 8'h00;
/*054*/LanguageConstructsTestSource_SOC_Array[84] = 8'h00;
/*055*/LanguageConstructsTestSource_SOC_Array[85] = 8'h00;
/*056*/LanguageConstructsTestSource_SOC_Array[86] = 8'h00;
/*057*/LanguageConstructsTestSource_SOC_Array[87] = 8'h00;
/*058*/LanguageConstructsTestSource_SOC_Array[88] = 8'h00;
/*059*/LanguageConstructsTestSource_SOC_Array[89] = 8'h00;
/*05A*/LanguageConstructsTestSource_SOC_Array[90] = 8'h00;
/*05B*/LanguageConstructsTestSource_SOC_Array[91] = 8'h00;
/*05C*/LanguageConstructsTestSource_SOC_Array[92] = 8'h00;
/*05D*/LanguageConstructsTestSource_SOC_Array[93] = 8'h00;
/*05E*/LanguageConstructsTestSource_SOC_Array[94] = 8'h00;
/*05F*/LanguageConstructsTestSource_SOC_Array[95] = 8'h00;
/*060*/LanguageConstructsTestSource_SOC_Array[96] = 8'h00;
/*061*/LanguageConstructsTestSource_SOC_Array[97] = 8'h00;
/*062*/LanguageConstructsTestSource_SOC_Array[98] = 8'h00;
/*063*/LanguageConstructsTestSource_SOC_Array[99] = 8'h00;
/*064*/LanguageConstructsTestSource_SOC_Array[100] = 8'h00;
/*065*/LanguageConstructsTestSource_SOC_Array[101] = 8'h00;
/*066*/LanguageConstructsTestSource_SOC_Array[102] = 8'h00;
/*067*/LanguageConstructsTestSource_SOC_Array[103] = 8'h00;
/*068*/LanguageConstructsTestSource_SOC_Array[104] = 8'h00;
/*069*/LanguageConstructsTestSource_SOC_Array[105] = 8'h00;
/*06A*/LanguageConstructsTestSource_SOC_Array[106] = 8'h00;
/*06B*/LanguageConstructsTestSource_SOC_Array[107] = 8'h00;
/*06C*/LanguageConstructsTestSource_SOC_Array[108] = 8'h00;
/*06D*/LanguageConstructsTestSource_SOC_Array[109] = 8'h00;
/*06E*/LanguageConstructsTestSource_SOC_Array[110] = 8'h00;
/*06F*/LanguageConstructsTestSource_SOC_Array[111] = 8'h00;
/*070*/LanguageConstructsTestSource_SOC_Array[112] = 8'h00;
/*071*/LanguageConstructsTestSource_SOC_Array[113] = 8'h00;
/*072*/LanguageConstructsTestSource_SOC_Array[114] = 8'h00;
/*073*/LanguageConstructsTestSource_SOC_Array[115] = 8'h00;
/*074*/LanguageConstructsTestSource_SOC_Array[116] = 8'h00;
/*075*/LanguageConstructsTestSource_SOC_Array[117] = 8'h00;
/*076*/LanguageConstructsTestSource_SOC_Array[118] = 8'h00;
/*077*/LanguageConstructsTestSource_SOC_Array[119] = 8'h00;
/*078*/LanguageConstructsTestSource_SOC_Array[120] = 8'h00;
/*079*/LanguageConstructsTestSource_SOC_Array[121] = 8'h00;
/*07A*/LanguageConstructsTestSource_SOC_Array[122] = 8'h00;
/*07B*/LanguageConstructsTestSource_SOC_Array[123] = 8'h00;
/*07C*/LanguageConstructsTestSource_SOC_Array[124] = 8'h00;
/*07D*/LanguageConstructsTestSource_SOC_Array[125] = 8'h00;
/*07E*/LanguageConstructsTestSource_SOC_Array[126] = 8'h00;
/*07F*/LanguageConstructsTestSource_SOC_Array[127] = 8'h00;
/*080*/LanguageConstructsTestSource_SOC_Array[128] = 8'h00;
/*081*/LanguageConstructsTestSource_SOC_Array[129] = 8'h00;
/*082*/LanguageConstructsTestSource_SOC_Array[130] = 8'h00;
/*083*/LanguageConstructsTestSource_SOC_Array[131] = 8'h00;
/*084*/LanguageConstructsTestSource_SOC_Array[132] = 8'h00;
/*085*/LanguageConstructsTestSource_SOC_Array[133] = 8'h00;
/*086*/LanguageConstructsTestSource_SOC_Array[134] = 8'h00;
/*087*/LanguageConstructsTestSource_SOC_Array[135] = 8'h00;
/*088*/LanguageConstructsTestSource_SOC_Array[136] = 8'h00;
/*089*/LanguageConstructsTestSource_SOC_Array[137] = 8'h00;
/*08A*/LanguageConstructsTestSource_SOC_Array[138] = 8'h00;
/*08B*/LanguageConstructsTestSource_SOC_Array[139] = 8'h00;
/*08C*/LanguageConstructsTestSource_SOC_Array[140] = 8'h00;
/*08D*/LanguageConstructsTestSource_SOC_Array[141] = 8'h00;
/*08E*/LanguageConstructsTestSource_SOC_Array[142] = 8'h00;
/*08F*/LanguageConstructsTestSource_SOC_Array[143] = 8'h00;
/*090*/LanguageConstructsTestSource_SOC_Array[144] = 8'h00;
/*091*/LanguageConstructsTestSource_SOC_Array[145] = 8'h00;
/*092*/LanguageConstructsTestSource_SOC_Array[146] = 8'h00;
/*093*/LanguageConstructsTestSource_SOC_Array[147] = 8'h00;
/*094*/LanguageConstructsTestSource_SOC_Array[148] = 8'h00;
/*095*/LanguageConstructsTestSource_SOC_Array[149] = 8'h00;
/*096*/LanguageConstructsTestSource_SOC_Array[150] = 8'h00;
/*097*/LanguageConstructsTestSource_SOC_Array[151] = 8'h00;
/*098*/LanguageConstructsTestSource_SOC_Array[152] = 8'h00;
/*099*/LanguageConstructsTestSource_SOC_Array[153] = 8'h00;
/*09A*/LanguageConstructsTestSource_SOC_Array[154] = 8'h00;
/*09B*/LanguageConstructsTestSource_SOC_Array[155] = 8'h00;
/*09C*/LanguageConstructsTestSource_SOC_Array[156] = 8'h00;
/*09D*/LanguageConstructsTestSource_SOC_Array[157] = 8'h00;
/*09E*/LanguageConstructsTestSource_SOC_Array[158] = 8'h00;
/*09F*/LanguageConstructsTestSource_SOC_Array[159] = 8'h00;
/*0A0*/LanguageConstructsTestSource_SOC_Array[160] = 8'h00;
/*0A1*/LanguageConstructsTestSource_SOC_Array[161] = 8'h00;
/*0A2*/LanguageConstructsTestSource_SOC_Array[162] = 8'h00;
/*0A3*/LanguageConstructsTestSource_SOC_Array[163] = 8'h00;
/*0A4*/LanguageConstructsTestSource_SOC_Array[164] = 8'h00;
/*0A5*/LanguageConstructsTestSource_SOC_Array[165] = 8'h00;
/*0A6*/LanguageConstructsTestSource_SOC_Array[166] = 8'h00;
/*0A7*/LanguageConstructsTestSource_SOC_Array[167] = 8'h00;
/*0A8*/LanguageConstructsTestSource_SOC_Array[168] = 8'h00;
/*0A9*/LanguageConstructsTestSource_SOC_Array[169] = 8'h00;
/*0AA*/LanguageConstructsTestSource_SOC_Array[170] = 8'h00;
/*0AB*/LanguageConstructsTestSource_SOC_Array[171] = 8'h00;
/*0AC*/LanguageConstructsTestSource_SOC_Array[172] = 8'h00;
/*0AD*/LanguageConstructsTestSource_SOC_Array[173] = 8'h00;
/*0AE*/LanguageConstructsTestSource_SOC_Array[174] = 8'h00;
/*0AF*/LanguageConstructsTestSource_SOC_Array[175] = 8'h00;
/*0B0*/LanguageConstructsTestSource_SOC_Array[176] = 8'h00;
/*0B1*/LanguageConstructsTestSource_SOC_Array[177] = 8'h00;
/*0B2*/LanguageConstructsTestSource_SOC_Array[178] = 8'h00;
/*0B3*/LanguageConstructsTestSource_SOC_Array[179] = 8'h00;
/*0B4*/LanguageConstructsTestSource_SOC_Array[180] = 8'h00;
/*0B5*/LanguageConstructsTestSource_SOC_Array[181] = 8'h00;
/*0B6*/LanguageConstructsTestSource_SOC_Array[182] = 8'h00;
/*0B7*/LanguageConstructsTestSource_SOC_Array[183] = 8'h00;
/*0B8*/LanguageConstructsTestSource_SOC_Array[184] = 8'h00;
/*0B9*/LanguageConstructsTestSource_SOC_Array[185] = 8'h00;
/*0BA*/LanguageConstructsTestSource_SOC_Array[186] = 8'h00;
/*0BB*/LanguageConstructsTestSource_SOC_Array[187] = 8'h00;
/*0BC*/LanguageConstructsTestSource_SOC_Array[188] = 8'h00;
/*0BD*/LanguageConstructsTestSource_SOC_Array[189] = 8'h00;
/*0BE*/LanguageConstructsTestSource_SOC_Array[190] = 8'h00;
/*0BF*/LanguageConstructsTestSource_SOC_Array[191] = 8'h00;
/*0C0*/LanguageConstructsTestSource_SOC_Array[192] = 8'h00;
/*0C1*/LanguageConstructsTestSource_SOC_Array[193] = 8'h00;
/*0C2*/LanguageConstructsTestSource_SOC_Array[194] = 8'h00;
/*0C3*/LanguageConstructsTestSource_SOC_Array[195] = 8'h00;
/*0C4*/LanguageConstructsTestSource_SOC_Array[196] = 8'h00;
/*0C5*/LanguageConstructsTestSource_SOC_Array[197] = 8'h00;
/*0C6*/LanguageConstructsTestSource_SOC_Array[198] = 8'h00;
/*0C7*/LanguageConstructsTestSource_SOC_Array[199] = 8'h00;
/*0C8*/LanguageConstructsTestSource_SOC_Array[200] = 8'h00;
/*0C9*/LanguageConstructsTestSource_SOC_Array[201] = 8'h00;
/*0CA*/LanguageConstructsTestSource_SOC_Array[202] = 8'h00;
/*0CB*/LanguageConstructsTestSource_SOC_Array[203] = 8'h00;
/*0CC*/LanguageConstructsTestSource_SOC_Array[204] = 8'h00;
/*0CD*/LanguageConstructsTestSource_SOC_Array[205] = 8'h00;
/*0CE*/LanguageConstructsTestSource_SOC_Array[206] = 8'h00;
/*0CF*/LanguageConstructsTestSource_SOC_Array[207] = 8'h00;
/*0D0*/LanguageConstructsTestSource_SOC_Array[208] = 8'h00;
/*0D1*/LanguageConstructsTestSource_SOC_Array[209] = 8'h00;
/*0D2*/LanguageConstructsTestSource_SOC_Array[210] = 8'h00;
/*0D3*/LanguageConstructsTestSource_SOC_Array[211] = 8'h00;
/*0D4*/LanguageConstructsTestSource_SOC_Array[212] = 8'h00;
/*0D5*/LanguageConstructsTestSource_SOC_Array[213] = 8'h00;
/*0D6*/LanguageConstructsTestSource_SOC_Array[214] = 8'h00;
/*0D7*/LanguageConstructsTestSource_SOC_Array[215] = 8'h00;
/*0D8*/LanguageConstructsTestSource_SOC_Array[216] = 8'h00;
/*0D9*/LanguageConstructsTestSource_SOC_Array[217] = 8'h00;
/*0DA*/LanguageConstructsTestSource_SOC_Array[218] = 8'h00;
/*0DB*/LanguageConstructsTestSource_SOC_Array[219] = 8'h00;
/*0DC*/LanguageConstructsTestSource_SOC_Array[220] = 8'h00;
/*0DD*/LanguageConstructsTestSource_SOC_Array[221] = 8'h00;
/*0DE*/LanguageConstructsTestSource_SOC_Array[222] = 8'h00;
/*0DF*/LanguageConstructsTestSource_SOC_Array[223] = 8'h00;
/*0E0*/LanguageConstructsTestSource_SOC_Array[224] = 8'h00;
/*0E1*/LanguageConstructsTestSource_SOC_Array[225] = 8'h00;
/*0E2*/LanguageConstructsTestSource_SOC_Array[226] = 8'h00;
/*0E3*/LanguageConstructsTestSource_SOC_Array[227] = 8'h00;
/*0E4*/LanguageConstructsTestSource_SOC_Array[228] = 8'h00;
/*0E5*/LanguageConstructsTestSource_SOC_Array[229] = 8'h00;
/*0E6*/LanguageConstructsTestSource_SOC_Array[230] = 8'h00;
/*0E7*/LanguageConstructsTestSource_SOC_Array[231] = 8'h00;
/*0E8*/LanguageConstructsTestSource_SOC_Array[232] = 8'h00;
/*0E9*/LanguageConstructsTestSource_SOC_Array[233] = 8'h00;
/*0EA*/LanguageConstructsTestSource_SOC_Array[234] = 8'h00;
/*0EB*/LanguageConstructsTestSource_SOC_Array[235] = 8'h00;
/*0EC*/LanguageConstructsTestSource_SOC_Array[236] = 8'h00;
/*0ED*/LanguageConstructsTestSource_SOC_Array[237] = 8'h00;
/*0EE*/LanguageConstructsTestSource_SOC_Array[238] = 8'h00;
/*0EF*/LanguageConstructsTestSource_SOC_Array[239] = 8'h00;
/*0F0*/LanguageConstructsTestSource_SOC_Array[240] = 8'h00;
/*0F1*/LanguageConstructsTestSource_SOC_Array[241] = 8'h00;
/*0F2*/LanguageConstructsTestSource_SOC_Array[242] = 8'h00;
/*0F3*/LanguageConstructsTestSource_SOC_Array[243] = 8'h00;
/*0F4*/LanguageConstructsTestSource_SOC_Array[244] = 8'h00;
/*0F5*/LanguageConstructsTestSource_SOC_Array[245] = 8'h00;
/*0F6*/LanguageConstructsTestSource_SOC_Array[246] = 8'h00;
/*0F7*/LanguageConstructsTestSource_SOC_Array[247] = 8'h00;
/*0F8*/LanguageConstructsTestSource_SOC_Array[248] = 8'h00;
/*0F9*/LanguageConstructsTestSource_SOC_Array[249] = 8'h00;
/*0FA*/LanguageConstructsTestSource_SOC_Array[250] = 8'h00;
/*0FB*/LanguageConstructsTestSource_SOC_Array[251] = 8'h00;
/*0FC*/LanguageConstructsTestSource_SOC_Array[252] = 8'h00;
/*0FD*/LanguageConstructsTestSource_SOC_Array[253] = 8'h00;
/*0FE*/LanguageConstructsTestSource_SOC_Array[254] = 8'h00;
/*0FF*/LanguageConstructsTestSource_SOC_Array[255] = 8'h00;
/*100*/LanguageConstructsTestSource_SOC_Array[256] = 8'h00;
/*101*/LanguageConstructsTestSource_SOC_Array[257] = 8'h00;
/*102*/LanguageConstructsTestSource_SOC_Array[258] = 8'h00;
/*103*/LanguageConstructsTestSource_SOC_Array[259] = 8'h00;
/*104*/LanguageConstructsTestSource_SOC_Array[260] = 8'h00;
/*105*/LanguageConstructsTestSource_SOC_Array[261] = 8'h00;
/*106*/LanguageConstructsTestSource_SOC_Array[262] = 8'h00;
/*107*/LanguageConstructsTestSource_SOC_Array[263] = 8'h00;
/*108*/LanguageConstructsTestSource_SOC_Array[264] = 8'h00;
/*109*/LanguageConstructsTestSource_SOC_Array[265] = 8'h00;
/*10A*/LanguageConstructsTestSource_SOC_Array[266] = 8'h00;
/*10B*/LanguageConstructsTestSource_SOC_Array[267] = 8'h00;
/*10C*/LanguageConstructsTestSource_SOC_Array[268] = 8'h00;
/*10D*/LanguageConstructsTestSource_SOC_Array[269] = 8'h00;
/*10E*/LanguageConstructsTestSource_SOC_Array[270] = 8'h00;
/*10F*/LanguageConstructsTestSource_SOC_Array[271] = 8'h00;
/*110*/LanguageConstructsTestSource_SOC_Array[272] = 8'h00;
/*111*/LanguageConstructsTestSource_SOC_Array[273] = 8'h00;
/*112*/LanguageConstructsTestSource_SOC_Array[274] = 8'h00;
/*113*/LanguageConstructsTestSource_SOC_Array[275] = 8'h00;
/*114*/LanguageConstructsTestSource_SOC_Array[276] = 8'h00;
/*115*/LanguageConstructsTestSource_SOC_Array[277] = 8'h00;
/*116*/LanguageConstructsTestSource_SOC_Array[278] = 8'h00;
/*117*/LanguageConstructsTestSource_SOC_Array[279] = 8'h00;
/*118*/LanguageConstructsTestSource_SOC_Array[280] = 8'h00;
/*119*/LanguageConstructsTestSource_SOC_Array[281] = 8'h00;
/*11A*/LanguageConstructsTestSource_SOC_Array[282] = 8'h00;
/*11B*/LanguageConstructsTestSource_SOC_Array[283] = 8'h00;
/*11C*/LanguageConstructsTestSource_SOC_Array[284] = 8'h00;
/*11D*/LanguageConstructsTestSource_SOC_Array[285] = 8'h00;
/*11E*/LanguageConstructsTestSource_SOC_Array[286] = 8'h00;
/*11F*/LanguageConstructsTestSource_SOC_Array[287] = 8'h00;
/*120*/LanguageConstructsTestSource_SOC_Array[288] = 8'h00;
/*121*/LanguageConstructsTestSource_SOC_Array[289] = 8'h00;
/*122*/LanguageConstructsTestSource_SOC_Array[290] = 8'h00;
/*123*/LanguageConstructsTestSource_SOC_Array[291] = 8'h00;
/*124*/LanguageConstructsTestSource_SOC_Array[292] = 8'h00;
/*125*/LanguageConstructsTestSource_SOC_Array[293] = 8'h00;
/*126*/LanguageConstructsTestSource_SOC_Array[294] = 8'h00;
/*127*/LanguageConstructsTestSource_SOC_Array[295] = 8'h00;
/*128*/LanguageConstructsTestSource_SOC_Array[296] = 8'h00;
/*129*/LanguageConstructsTestSource_SOC_Array[297] = 8'h00;
/*12A*/LanguageConstructsTestSource_SOC_Array[298] = 8'h00;
/*12B*/LanguageConstructsTestSource_SOC_Array[299] = 8'h00;
/*12C*/LanguageConstructsTestSource_SOC_Array[300] = 8'h00;
/*12D*/LanguageConstructsTestSource_SOC_Array[301] = 8'h00;
/*12E*/LanguageConstructsTestSource_SOC_Array[302] = 8'h00;
/*12F*/LanguageConstructsTestSource_SOC_Array[303] = 8'h00;
/*130*/LanguageConstructsTestSource_SOC_Array[304] = 8'h00;
/*131*/LanguageConstructsTestSource_SOC_Array[305] = 8'h00;
/*132*/LanguageConstructsTestSource_SOC_Array[306] = 8'h00;
/*133*/LanguageConstructsTestSource_SOC_Array[307] = 8'h00;
/*134*/LanguageConstructsTestSource_SOC_Array[308] = 8'h00;
/*135*/LanguageConstructsTestSource_SOC_Array[309] = 8'h00;
/*136*/LanguageConstructsTestSource_SOC_Array[310] = 8'h00;
/*137*/LanguageConstructsTestSource_SOC_Array[311] = 8'h00;
/*138*/LanguageConstructsTestSource_SOC_Array[312] = 8'h00;
/*139*/LanguageConstructsTestSource_SOC_Array[313] = 8'h00;
/*13A*/LanguageConstructsTestSource_SOC_Array[314] = 8'h00;
/*13B*/LanguageConstructsTestSource_SOC_Array[315] = 8'h00;
/*13C*/LanguageConstructsTestSource_SOC_Array[316] = 8'h00;
/*13D*/LanguageConstructsTestSource_SOC_Array[317] = 8'h00;
/*13E*/LanguageConstructsTestSource_SOC_Array[318] = 8'h00;
/*13F*/LanguageConstructsTestSource_SOC_Array[319] = 8'h00;
/*140*/LanguageConstructsTestSource_SOC_Array[320] = 8'h00;
/*141*/LanguageConstructsTestSource_SOC_Array[321] = 8'h00;
/*142*/LanguageConstructsTestSource_SOC_Array[322] = 8'h00;
/*143*/LanguageConstructsTestSource_SOC_Array[323] = 8'h00;
/*144*/LanguageConstructsTestSource_SOC_Array[324] = 8'h00;
/*145*/LanguageConstructsTestSource_SOC_Array[325] = 8'h00;
/*146*/LanguageConstructsTestSource_SOC_Array[326] = 8'h00;
/*147*/LanguageConstructsTestSource_SOC_Array[327] = 8'h00;
/*148*/LanguageConstructsTestSource_SOC_Array[328] = 8'h00;
/*149*/LanguageConstructsTestSource_SOC_Array[329] = 8'h00;
/*14A*/LanguageConstructsTestSource_SOC_Array[330] = 8'h00;
/*14B*/LanguageConstructsTestSource_SOC_Array[331] = 8'h00;
/*14C*/LanguageConstructsTestSource_SOC_Array[332] = 8'h00;
/*14D*/LanguageConstructsTestSource_SOC_Array[333] = 8'h00;
/*14E*/LanguageConstructsTestSource_SOC_Array[334] = 8'h00;
/*14F*/LanguageConstructsTestSource_SOC_Array[335] = 8'h00;
/*150*/LanguageConstructsTestSource_SOC_Array[336] = 8'h00;
/*151*/LanguageConstructsTestSource_SOC_Array[337] = 8'h00;
/*152*/LanguageConstructsTestSource_SOC_Array[338] = 8'h00;
/*153*/LanguageConstructsTestSource_SOC_Array[339] = 8'h00;
/*154*/LanguageConstructsTestSource_SOC_Array[340] = 8'h00;
/*155*/LanguageConstructsTestSource_SOC_Array[341] = 8'h00;
/*156*/LanguageConstructsTestSource_SOC_Array[342] = 8'h00;
/*157*/LanguageConstructsTestSource_SOC_Array[343] = 8'h00;
/*158*/LanguageConstructsTestSource_SOC_Array[344] = 8'h00;
/*159*/LanguageConstructsTestSource_SOC_Array[345] = 8'h00;
/*15A*/LanguageConstructsTestSource_SOC_Array[346] = 8'h00;
/*15B*/LanguageConstructsTestSource_SOC_Array[347] = 8'h00;
/*15C*/LanguageConstructsTestSource_SOC_Array[348] = 8'h00;
/*15D*/LanguageConstructsTestSource_SOC_Array[349] = 8'h00;
/*15E*/LanguageConstructsTestSource_SOC_Array[350] = 8'h00;
/*15F*/LanguageConstructsTestSource_SOC_Array[351] = 8'h00;
/*160*/LanguageConstructsTestSource_SOC_Array[352] = 8'h00;
/*161*/LanguageConstructsTestSource_SOC_Array[353] = 8'h00;
/*162*/LanguageConstructsTestSource_SOC_Array[354] = 8'h00;
/*163*/LanguageConstructsTestSource_SOC_Array[355] = 8'h00;
/*164*/LanguageConstructsTestSource_SOC_Array[356] = 8'h00;
/*165*/LanguageConstructsTestSource_SOC_Array[357] = 8'h00;
/*166*/LanguageConstructsTestSource_SOC_Array[358] = 8'h00;
/*167*/LanguageConstructsTestSource_SOC_Array[359] = 8'h00;
/*168*/LanguageConstructsTestSource_SOC_Array[360] = 8'h00;
/*169*/LanguageConstructsTestSource_SOC_Array[361] = 8'h00;
/*16A*/LanguageConstructsTestSource_SOC_Array[362] = 8'h00;
/*16B*/LanguageConstructsTestSource_SOC_Array[363] = 8'h00;
/*16C*/LanguageConstructsTestSource_SOC_Array[364] = 8'h00;
/*16D*/LanguageConstructsTestSource_SOC_Array[365] = 8'h00;
/*16E*/LanguageConstructsTestSource_SOC_Array[366] = 8'h00;
/*16F*/LanguageConstructsTestSource_SOC_Array[367] = 8'h00;
/*170*/LanguageConstructsTestSource_SOC_Array[368] = 8'h00;
/*171*/LanguageConstructsTestSource_SOC_Array[369] = 8'h00;
/*172*/LanguageConstructsTestSource_SOC_Array[370] = 8'h00;
/*173*/LanguageConstructsTestSource_SOC_Array[371] = 8'h00;
/*174*/LanguageConstructsTestSource_SOC_Array[372] = 8'h00;
/*175*/LanguageConstructsTestSource_SOC_Array[373] = 8'h00;
/*176*/LanguageConstructsTestSource_SOC_Array[374] = 8'h00;
/*177*/LanguageConstructsTestSource_SOC_Array[375] = 8'h00;
/*178*/LanguageConstructsTestSource_SOC_Array[376] = 8'h00;
/*179*/LanguageConstructsTestSource_SOC_Array[377] = 8'h00;
/*17A*/LanguageConstructsTestSource_SOC_Array[378] = 8'h00;
/*17B*/LanguageConstructsTestSource_SOC_Array[379] = 8'h00;
/*17C*/LanguageConstructsTestSource_SOC_Array[380] = 8'h00;
/*17D*/LanguageConstructsTestSource_SOC_Array[381] = 8'h00;
/*17E*/LanguageConstructsTestSource_SOC_Array[382] = 8'h00;
/*17F*/LanguageConstructsTestSource_SOC_Array[383] = 8'h00;
/*180*/LanguageConstructsTestSource_SOC_Array[384] = 8'h00;
/*181*/LanguageConstructsTestSource_SOC_Array[385] = 8'h00;
/*182*/LanguageConstructsTestSource_SOC_Array[386] = 8'h00;
/*183*/LanguageConstructsTestSource_SOC_Array[387] = 8'h00;
/*184*/LanguageConstructsTestSource_SOC_Array[388] = 8'h00;
/*185*/LanguageConstructsTestSource_SOC_Array[389] = 8'h00;
/*186*/LanguageConstructsTestSource_SOC_Array[390] = 8'h00;
/*187*/LanguageConstructsTestSource_SOC_Array[391] = 8'h00;
/*188*/LanguageConstructsTestSource_SOC_Array[392] = 8'h00;
/*189*/LanguageConstructsTestSource_SOC_Array[393] = 8'h00;
/*18A*/LanguageConstructsTestSource_SOC_Array[394] = 8'h00;
/*18B*/LanguageConstructsTestSource_SOC_Array[395] = 8'h00;
/*18C*/LanguageConstructsTestSource_SOC_Array[396] = 8'h00;
/*18D*/LanguageConstructsTestSource_SOC_Array[397] = 8'h00;
/*18E*/LanguageConstructsTestSource_SOC_Array[398] = 8'h00;
/*18F*/LanguageConstructsTestSource_SOC_Array[399] = 8'h00;
/*190*/LanguageConstructsTestSource_SOC_Array[400] = 8'h00;
/*191*/LanguageConstructsTestSource_SOC_Array[401] = 8'h00;
/*192*/LanguageConstructsTestSource_SOC_Array[402] = 8'h00;
/*193*/LanguageConstructsTestSource_SOC_Array[403] = 8'h00;
/*194*/LanguageConstructsTestSource_SOC_Array[404] = 8'h00;
/*195*/LanguageConstructsTestSource_SOC_Array[405] = 8'h00;
/*196*/LanguageConstructsTestSource_SOC_Array[406] = 8'h00;
/*197*/LanguageConstructsTestSource_SOC_Array[407] = 8'h00;
/*198*/LanguageConstructsTestSource_SOC_Array[408] = 8'h00;
/*199*/LanguageConstructsTestSource_SOC_Array[409] = 8'h00;
/*19A*/LanguageConstructsTestSource_SOC_Array[410] = 8'h00;
/*19B*/LanguageConstructsTestSource_SOC_Array[411] = 8'h00;
/*19C*/LanguageConstructsTestSource_SOC_Array[412] = 8'h00;
/*19D*/LanguageConstructsTestSource_SOC_Array[413] = 8'h00;
/*19E*/LanguageConstructsTestSource_SOC_Array[414] = 8'h00;
/*19F*/LanguageConstructsTestSource_SOC_Array[415] = 8'h00;
/*1A0*/LanguageConstructsTestSource_SOC_Array[416] = 8'h00;
/*1A1*/LanguageConstructsTestSource_SOC_Array[417] = 8'h00;
/*1A2*/LanguageConstructsTestSource_SOC_Array[418] = 8'h00;
/*1A3*/LanguageConstructsTestSource_SOC_Array[419] = 8'h00;
/*1A4*/LanguageConstructsTestSource_SOC_Array[420] = 8'h00;
/*1A5*/LanguageConstructsTestSource_SOC_Array[421] = 8'h00;
/*1A6*/LanguageConstructsTestSource_SOC_Array[422] = 8'h00;
/*1A7*/LanguageConstructsTestSource_SOC_Array[423] = 8'h00;
/*1A8*/LanguageConstructsTestSource_SOC_Array[424] = 8'h00;
/*1A9*/LanguageConstructsTestSource_SOC_Array[425] = 8'h00;
/*1AA*/LanguageConstructsTestSource_SOC_Array[426] = 8'h00;
/*1AB*/LanguageConstructsTestSource_SOC_Array[427] = 8'h00;
/*1AC*/LanguageConstructsTestSource_SOC_Array[428] = 8'h00;
/*1AD*/LanguageConstructsTestSource_SOC_Array[429] = 8'h00;
/*1AE*/LanguageConstructsTestSource_SOC_Array[430] = 8'h00;
/*1AF*/LanguageConstructsTestSource_SOC_Array[431] = 8'h00;
/*1B0*/LanguageConstructsTestSource_SOC_Array[432] = 8'h00;
/*1B1*/LanguageConstructsTestSource_SOC_Array[433] = 8'h00;
/*1B2*/LanguageConstructsTestSource_SOC_Array[434] = 8'h00;
/*1B3*/LanguageConstructsTestSource_SOC_Array[435] = 8'h00;
/*1B4*/LanguageConstructsTestSource_SOC_Array[436] = 8'h00;
/*1B5*/LanguageConstructsTestSource_SOC_Array[437] = 8'h00;
/*1B6*/LanguageConstructsTestSource_SOC_Array[438] = 8'h00;
/*1B7*/LanguageConstructsTestSource_SOC_Array[439] = 8'h00;
/*1B8*/LanguageConstructsTestSource_SOC_Array[440] = 8'h00;
/*1B9*/LanguageConstructsTestSource_SOC_Array[441] = 8'h00;
/*1BA*/LanguageConstructsTestSource_SOC_Array[442] = 8'h00;
/*1BB*/LanguageConstructsTestSource_SOC_Array[443] = 8'h00;
/*1BC*/LanguageConstructsTestSource_SOC_Array[444] = 8'h00;
/*1BD*/LanguageConstructsTestSource_SOC_Array[445] = 8'h00;
/*1BE*/LanguageConstructsTestSource_SOC_Array[446] = 8'h00;
/*1BF*/LanguageConstructsTestSource_SOC_Array[447] = 8'h00;
/*1C0*/LanguageConstructsTestSource_SOC_Array[448] = 8'h00;
/*1C1*/LanguageConstructsTestSource_SOC_Array[449] = 8'h00;
/*1C2*/LanguageConstructsTestSource_SOC_Array[450] = 8'h00;
/*1C3*/LanguageConstructsTestSource_SOC_Array[451] = 8'h00;
/*1C4*/LanguageConstructsTestSource_SOC_Array[452] = 8'h00;
/*1C5*/LanguageConstructsTestSource_SOC_Array[453] = 8'h00;
/*1C6*/LanguageConstructsTestSource_SOC_Array[454] = 8'h00;
/*1C7*/LanguageConstructsTestSource_SOC_Array[455] = 8'h00;
/*1C8*/LanguageConstructsTestSource_SOC_Array[456] = 8'h00;
/*1C9*/LanguageConstructsTestSource_SOC_Array[457] = 8'h00;
/*1CA*/LanguageConstructsTestSource_SOC_Array[458] = 8'h00;
/*1CB*/LanguageConstructsTestSource_SOC_Array[459] = 8'h00;
/*1CC*/LanguageConstructsTestSource_SOC_Array[460] = 8'h00;
/*1CD*/LanguageConstructsTestSource_SOC_Array[461] = 8'h00;
/*1CE*/LanguageConstructsTestSource_SOC_Array[462] = 8'h00;
/*1CF*/LanguageConstructsTestSource_SOC_Array[463] = 8'h00;
/*1D0*/LanguageConstructsTestSource_SOC_Array[464] = 8'h00;
/*1D1*/LanguageConstructsTestSource_SOC_Array[465] = 8'h00;
/*1D2*/LanguageConstructsTestSource_SOC_Array[466] = 8'h00;
/*1D3*/LanguageConstructsTestSource_SOC_Array[467] = 8'h00;
/*1D4*/LanguageConstructsTestSource_SOC_Array[468] = 8'h00;
/*1D5*/LanguageConstructsTestSource_SOC_Array[469] = 8'h00;
/*1D6*/LanguageConstructsTestSource_SOC_Array[470] = 8'h00;
/*1D7*/LanguageConstructsTestSource_SOC_Array[471] = 8'h00;
/*1D8*/LanguageConstructsTestSource_SOC_Array[472] = 8'h00;
/*1D9*/LanguageConstructsTestSource_SOC_Array[473] = 8'h00;
/*1DA*/LanguageConstructsTestSource_SOC_Array[474] = 8'h00;
/*1DB*/LanguageConstructsTestSource_SOC_Array[475] = 8'h00;
/*1DC*/LanguageConstructsTestSource_SOC_Array[476] = 8'h00;
/*1DD*/LanguageConstructsTestSource_SOC_Array[477] = 8'h00;
/*1DE*/LanguageConstructsTestSource_SOC_Array[478] = 8'h00;
/*1DF*/LanguageConstructsTestSource_SOC_Array[479] = 8'h00;
/*1E0*/LanguageConstructsTestSource_SOC_Array[480] = 8'h00;
/*1E1*/LanguageConstructsTestSource_SOC_Array[481] = 8'h00;
/*1E2*/LanguageConstructsTestSource_SOC_Array[482] = 8'h00;
/*1E3*/LanguageConstructsTestSource_SOC_Array[483] = 8'h00;
/*1E4*/LanguageConstructsTestSource_SOC_Array[484] = 8'h00;
/*1E5*/LanguageConstructsTestSource_SOC_Array[485] = 8'h00;
/*1E6*/LanguageConstructsTestSource_SOC_Array[486] = 8'h00;
/*1E7*/LanguageConstructsTestSource_SOC_Array[487] = 8'h00;
/*1E8*/LanguageConstructsTestSource_SOC_Array[488] = 8'h00;
/*1E9*/LanguageConstructsTestSource_SOC_Array[489] = 8'h00;
/*1EA*/LanguageConstructsTestSource_SOC_Array[490] = 8'h00;
/*1EB*/LanguageConstructsTestSource_SOC_Array[491] = 8'h00;
/*1EC*/LanguageConstructsTestSource_SOC_Array[492] = 8'h00;
/*1ED*/LanguageConstructsTestSource_SOC_Array[493] = 8'h00;
/*1EE*/LanguageConstructsTestSource_SOC_Array[494] = 8'h00;
/*1EF*/LanguageConstructsTestSource_SOC_Array[495] = 8'h00;
/*1F0*/LanguageConstructsTestSource_SOC_Array[496] = 8'h00;
/*1F1*/LanguageConstructsTestSource_SOC_Array[497] = 8'h00;
/*1F2*/LanguageConstructsTestSource_SOC_Array[498] = 8'h00;
/*1F3*/LanguageConstructsTestSource_SOC_Array[499] = 8'h00;
/*1F4*/LanguageConstructsTestSource_SOC_Array[500] = 8'h00;
/*1F5*/LanguageConstructsTestSource_SOC_Array[501] = 8'h00;
/*1F6*/LanguageConstructsTestSource_SOC_Array[502] = 8'h00;
/*1F7*/LanguageConstructsTestSource_SOC_Array[503] = 8'h00;
/*1F8*/LanguageConstructsTestSource_SOC_Array[504] = 8'h00;
/*1F9*/LanguageConstructsTestSource_SOC_Array[505] = 8'h00;
/*1FA*/LanguageConstructsTestSource_SOC_Array[506] = 8'h00;
/*1FB*/LanguageConstructsTestSource_SOC_Array[507] = 8'h00;
/*1FC*/LanguageConstructsTestSource_SOC_Array[508] = 8'h00;
/*1FD*/LanguageConstructsTestSource_SOC_Array[509] = 8'h00;
/*1FE*/LanguageConstructsTestSource_SOC_Array[510] = 8'h00;
/*1FF*/LanguageConstructsTestSource_SOC_Array[511] = 8'h00;

// END MEM_INIT
end

	
endmodule